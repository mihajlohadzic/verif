`ifndef CONFIGURATION_PKG_SV
 `define CONFIGURATION_PKG_SV

package configurations_pkg;
   import uvm_pkg::*;
 `include "uvm_macros.svh"
 `include "config.sv"
endpackage: configurations_pkg


`endif
